library ieee;
use ieee.std_logic_1164.all;

entity testbench3 is
end testbench3;

architecture tb of testbench3 is
	component watch
		port( reset, en, clk: in std_logic;
	y2,y1,y0: out std_logic_vector(3 downto 0));
	end component;
signal reset, en, clk: std_logic;
signal y2,y1,y0: std_logic_vector(3 downto 0);
begin 
	DUT: watch port map(reset, en, clk, y2, y1, y0);
	 process
		 begin
		 clk <= '0';
		 wait for 5 ns;
		 clk <= '1';
		 wait for 5 ns;
	 end process;
	 
	 process
		 begin
		 reset <= '1';
		 wait for 2 ns;
		 reset <= '0';
		 wait for 400 ns;
	 end process;
	 
	 process
		 begin
		 en <= '0';
		 wait for 5 ns;
		 en <= '1';
		 wait for 20 ns;
	 end process;
	
 end tb;